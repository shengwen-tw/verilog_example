`timescale 1ms/10us

module test_dff();
endmodule
